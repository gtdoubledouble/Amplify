CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
31 91 1244 738
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
31 91 1244 738
144179218 0
0
6 Title:
5 Name:
0
0
0
7
9 V Source~
197 154 185 0 1 5
0 0
0
0 0 17248 90
10 2.55V  Max
-35 -20 35 -12
3 PWM
-11 -30 10 -22
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
8953 0 0
0
0
7 Ground~
168 278 216 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
9 Resistor~
219 208 185 0 1 5
0 0
0
0 0 864 0
3 100
-10 -14 11 -6
1 R
-4 -24 3 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
9 Resistor~
219 278 121 0 1 5
0 0
0
0 0 8928 90
3 100
5 0 26 8
1 R
11 -10 18 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
4 LED~
171 278 155 0 1 2
10 0
0
0 0 368 0
9 LED STRIP
18 -4 81 4
0
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 0 0 0 0
1 D
5394 0 0
0
0
12 NPN Trans:C~
219 273 185 0 1 7
0 0
0
0 0 832 0
6 2N3904
17 0 59 8
3 NPN
27 -11 48 -3
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 0 0 0 0
1 Q
7734 0 0
0
0
2 +V
167 279 77 0 1 3
0 0
0
0 0 54240 0
3 12V
-10 -22 11 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
6
2 1 0 0 0 0 0 1 3 0 0 2
175 185
190 185
1 3 0 0 0 0 0 2 6 0 0 2
278 210
278 203
2 2 0 0 0 0 0 3 6 0 0 2
226 185
255 185
2 1 0 0 0 0 0 5 6 0 0 2
278 165
278 167
2 1 0 0 0 0 0 4 7 0 0 4
278 103
278 105
279 105
279 86
1 1 0 0 0 0 0 4 5 0 0 2
278 139
278 145
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
